
/*
 * Module 'cpu'
 *
 * Main module for kore-v
 */
module cpu;
  /* Define registers. */
  logic [31:0] pc;

  /* Define the regfile module. */

endmodule
