
/*
 * Module 'cpu'
 *
 * Main module for kore-v
 */
module cpu;
  /* Define registers. */
  logic [31:0] regfile[32];
  logic [31:0] pc;

endmodule
